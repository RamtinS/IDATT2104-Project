
module add(
    input [7:0] A, B,
    output [8:0] C
);

    assign C = A + B;
endmodule

